
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity hazard_detector is
    port (
        a : in std_logic_vector(31 downto 0)
    );
end hazard_detector;

architecture hazard_detector_arch of hazard_detector is

begin
end hazard_detector_arch;

